module server

import io
import net
import x.json2 as jsn
import src.db_utils as db

pub struct MessagramServer
{
	pub mut:
		host			string
		port 			int = 666

		clients			[]Client
		main_socket 	net.TcpListener
}

pub fn start_messagram_server(mut m MessagramServer)
{
	m.main_socket = net.listen_tcp(.ip6, ":${m.port}") or {
		println("[ X ], Error, Unable to start server....!")
		return
	}

	println("[ + ] Messagram server has been started....!")

	m.client_listener()
}

pub fn (mut m MessagramServer) client_listener() 
{
	for {
		mut client := m.main_socket.accept() or { &net.TcpConn{} }

		/*
		 	API LOGIN AUTHENICATION SHOULD ONLY COME FROM A SPECIFIC IP OR LOCALHOST
			IT WILL BE SENT TO PARSE AND AUTHORIZATION CHECKING 
		*/
		user_ip := client.peer_ip() or { "" }
		if user_ip == "BACKEND_IP_HERE" {
			m.authenicate_user(mut client)
		}
		m.client_authenticator(mut client)
	}
}

pub fn (mut m MessagramServer) authenicate_user(mut c net.TcpConn)
{
	mut reader := io.new_buffered_reader(reader: c)
	mut info := reader.read_line() or { "" }

	if !info.starts_with("{") && !info.ends_with("}") {
		// FORM A JSON RESPONSE
	}


}

/*
	A sessionID must be generated by authenicating via API Auth Endpoint
*/
pub fn (mut m MessagramServer) client_authenticator(mut c net.TcpConn) 
{
	mut reader := io.new_buffered_reader(reader: c)

	c.write_string("[ + ] Welcome to Messagram Server v0.0.1\n") or { 0 }
	login := reader.read_line() or { "" }

	println(login)
	if !login.starts_with("{") && !login.ends_with("}") {
		println("[ X ] Error, Invalid login data provided....!\r\n\t=> Disconnecting user " + c.peer_ip() or { "" } + "\r\n\t=>\r\n${login}")
		c.close() or { net.TcpConn{} }
		return 
	}

	/*	
		{

			"username": "",
			"password": "",
			"ip": "",
			"sid": ""
		}
	*/
	mut login_data := (jsn.raw_decode("${login}") or { jsn.Any{} }).as_map()

	if "cmd" !in login_data || "username" !in login_data || "sessionID" !in login_data || "hwid" !in login_data {
		println("[ X ] Error, Invalid JSON Response")
		c.close() or { net.TcpConn{} }
		return
	}

	cmd 		:= login_data['cmd'] or { "N/A" }
	username 	:= login_data['username'] or { "N/A" }
	sessionID	:= login_data['sessionID'] or { "N/A" }
	hwid 		:= login_data['hwid'] or { "N/A" }

	println("${username} ${password} ${ip} ${sid}")

	// Login Authenication
}

pub fn (mut m MessagramServer) command_handler(login_data string) 
{

}

/*
	[@DOC]
	pub fn (mut m MessagramServer) add_session_key(sid string, username string) string

	Generate a sessionID to return to user via API req to connect through a client
*/
pub fn (mut m MessagramServer) add_session_key(sid string, username string) string
{
	// find user profile 
	// generate a key to return 
	// add sessionid to profile 
	// append the profile to the MessagramServer struck
	// wait for 60 seconds before terminating the sessionID 
}