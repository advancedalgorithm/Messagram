module server

import io
import net
import time
import x.json2 as jsn

import src.db_utils as db

pub struct MessagramServer
{
	pub mut:
		host			string
		port 			int = 666
		users			[]db.User
		clients			[]Client
		main_socket 	net.TcpListener
}

pub fn start_messagram_server(mut m MessagramServer, mut users []db.User)
{
	m.main_socket = net.listen_tcp(.ip6, ":${m.port}") or {
		println("[ X ] Error, Unable to start server....!")
		return
	}

	m.users = users

	println("[ + ] Messagram server has been started....!")

	m.client_listener()
}

pub fn (mut m MessagramServer) client_listener() 
{
	for {
		mut client := m.main_socket.accept() or { &net.TcpConn{} }

		/*
		 	API LOGIN AUTHENICATION SHOULD ONLY COME FROM A SPECIFIC IP OR LOCALHOST
			IT WILL BE SENT TO PARSE AND AUTHORIZATION CHECKING 
		*/
		user_ip := client.peer_ip() or { "" }
		client.set_read_timeout(time.infinite)
		if user_ip == "BACKEND_IP_HERE" { // WEBSITE
			m.authenticate_user(mut client)
		}
		m.client_authenticator(mut client)
	}
}

/*
* USE FOR API ENDPOINT
*
* Authorize user then generate a sessionID for user on the API Endpoint
*
*/
pub fn (mut m MessagramServer) authenticate_user(mut c net.TcpConn)
{
	mut reader := io.new_buffered_reader(reader: c)
	mut info := reader.read_line() or { "" }

	if !info.starts_with("{") && !info.ends_with("}") {
		// FORM A JSON RESPONSE
	}


	// Find user
	// mut user, chk := authorize_user(username, password)

	// mut socket_client := new_client(mut c, 
	// m.clients << socket_client
}

/*
	A sessionID must be generated by authenicating via API Auth Endpoint
*/
pub fn (mut m MessagramServer) client_authenticator(mut c net.TcpConn) 
{
	mut reader := io.new_buffered_reader(reader: c)

	// c.write_string("[ + ] Welcome to Messagram Server v0.0.1\n") or { 0 }
	login := reader.read_line() or { "" }

	if !login.starts_with("{") && !login.ends_with("}") {
		println("[ X ] Error, Invalid login data provided....!\r\n\t=> Disconnecting user " + c.peer_ip() or { "" } + "\r\n\t=>\r\n${login}")
		c.close() or { return }
		return 
	}

	/*
		{
			"cmd_t": ""
			"username": "",
			"sid": "",
			"hwid": "",
			"client_name": "",
			"client_version": ""
		}
	*/
	mut login_data := (jsn.raw_decode("${login}") or { jsn.Any{} }).as_map()

	if "cmd_t" !in login_data || "username" !in login_data || "sid" !in login_data || "hwid" !in login_data {
		println("[ X ] Error, Invalid JSON Response")
		c.close() or { return }
		return
	}

	cmd 		:= (login_data['cmd_t'] 			or { "" }).str()
	username 	:= (login_data['username'] 			or { "" }).str()
	sid 		:= (login_data['sid'] 				or { "" }).str()
	hwid		:= (login_data['hwid'] 				or { "" }).str()
	client_name := (login_data['client_name']		or { "" }).str()
	client_v 	:= (login_data['client_version'] 	or { "" }).str()
	host_addr	:= c.peer_ip() or { "" }

	// Login Authenication
	mut user 		:= m.find_account(username)
	mut client, chk := m.find_client_id(sid, hwid)

	println(login_data)
	mut r := parse_cmd(mut client.info, login)
	mut new_resp := r.parse_cmd_data()

	println("Inbound Command: ${r.to_str()}")
	println("Outbound Command: ${new_resp.to_str()}")

	if !chk {
		c.write_string("{\"status\": \"false\", \"resp_t\": \"user_resp\", \"cmd_t\": \"INVALID_LOGIN_INFO\"}") or { 0 }
		c.close() or { return }
		return
	}

	/* Updating the Client's Socket && Client Information */
	client.socket 		= c
	client.using_app 	= true
	client.app_name 	= client_name
	client.app_version 	= client_v

	c.write_string("{\"status\": \"true\", \"resp_t\": \"user_resp\", \"cmd_t\": \"SUCCESSFUL_LOGIN\"}") or { 0 }
	m.command_handler(mut c, mut client)
}

/*
	Client Cmd Handler

	Handling account actions such as setting editing, dm actions etc
*/
pub fn (mut m MessagramServer) command_handler(mut socket net.TcpConn, mut client Client)
{
	mut reader := io.new_buffered_reader(reader: socket)
	for
	{
		new_data := reader.read_line() or {
			m.disconnect_user(mut client.socket)
			println("[ X ] Error, Client disconnected from socket\r\n\t=>${client.info.username}.....!")
			return
		}

		if !new_data.starts_with("{") || !new_data.ends_with("}")
		{
			m.disconnect_user(mut client.socket)
			println("[ X ] Error, Invalid JSON Data Received!")
			return
		}

		/*
			Default JSON Fields

			There will be additional keys to parse depending on the
			type of commands received
			{
				"cmd": "",
				"username": "",
				"sessionID": "",
				"hwid": "",
				"client_name": "",
				"client_version": ""
			}

			Validate the information below to check the connection
		*/
		json_data 	:= (jsn.raw_decode(new_data) 	or { jsn.Any{} }).as_map()
		cmd 		:= (json_data['cmd_t'] 			or { "" }).str()
		username 	:= (json_data['username'] 		or { "" }).str()
		sid 		:= (json_data['sessionID'] 		or { "" }).str()
		hwid 		:= (json_data['hwid'] 			or { "" }).str() 
		client_name	:= (json_data['client_name']	or { "" }).str()
		client_v	:= (json_data['client_v']		or { "" }).str() 

		// DO ALL CONNECTION VALIDATION CHECKS HERE

		mut r := parse_cmd(mut client.info, new_data)
		mut new_r := r.parse_cmd_data()


		println("Inbound Command: ${r.to_str()}")
		println("Outbound Command: ${new_r.to_str()}")

		/* UNCOMMENT THE FUNCTION BELOW ONCE ALL RESPONSES ARE FINISHED */
		
		// handle_command(mut socket, mut new_r)
		// socket.write_string("${new_r.to_str()}") or { 0 }
	}
}

pub fn (mut m MessagramServer) disconnect_user(mut socket net.TcpConn) bool
{
	socket.close() or { return false }

	for i, client in m.clients 
	{
		if client.socket == socket { m.clients.delete(i) }
	}

	return true
}

/*
	Find the client id in the (CONNECTED SOCKET CLIENTS) using sid

	Args:
		- sid: sessionID
	
	Returns:
		- Client structure
*/
pub fn (mut m MessagramServer) find_client_id(sid string, h string) (Client, bool)
{
	mut new := Client{socket: &net.TcpConn{}}
	for mut client in m.clients 
	{
		if client.sid == sid && client.hwid == h { return client, true }
	}

	return new, false
}

/* 
	Find an account within Messagram's Database (NOT CONNECTED SOCKET CLIENTS)
	
	Args:
		- username: string
	
	Returns:
		- User structure
*/
pub fn (mut m MessagramServer) find_account(username string) db.User
{
	println("Searching... ${username}")
	for mut user in m.users
	{
		if user.username == username { return user }
	}

	return db.User{}
}