module db_utils

pub const (
	user_dbpath = "assets/db/users.mg"
)