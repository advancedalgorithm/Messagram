module db_utils

pub struct Dm 
{
	pub mut:
		name		string
		user_id		string
		messages 	[]string
		
}