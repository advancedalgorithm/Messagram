module server

import os
import io
import net
import time
import x.json2 as jsn

import src.db_utils as db

pub struct MessagramServer
{
	pub mut:
		host			string
		port 			int = 666
		users			[]db.User
		clients			[]Client
		client_sockets  []net.TcpConn
		main_socket 	net.TcpListener
}

pub fn start_messagram_server(mut m MessagramServer, mut users []db.User)
{
	m.main_socket = net.listen_tcp(.ip6, ":${m.port}") or {
		println("[ X ] Error, Unable to start server....!")
		return
	}

	m.users = users

	println("[ + ] Messagram server has been started....!")

	m.client_listener()
}

pub fn (mut m MessagramServer) client_listener() 
{
	for {
		mut client := m.main_socket.accept() or { 
			println("[ X ] Unable to accept connection")
			return
		}

		/*
		 	API LOGIN AUTHENICATION SHOULD ONLY COME FROM A SPECIFIC IP OR LOCALHOST
			IT WILL BE SENT TO PARSE AND AUTHORIZATION CHECKING 
		*/
		user_ip := client.peer_ip() or { "" }
		client.set_read_timeout(time.infinite)
		if user_ip == "BACKEND_IP_HERE" { // WEBSITE
			spawn m.authenticate_user(mut client)
		}
		spawn m.client_authenticator(mut client)
	}
}

/*
* USE FOR API ENDPOINT
*
* Authorize user then generate a sessionID for user on the API Endpoint
*
*/
pub fn (mut m MessagramServer) authenticate_user(mut c net.TcpConn)
{
	mut reader := io.new_buffered_reader(reader: c)
	mut info := reader.read_line() or { "" }

	if !info.starts_with("{") && !info.ends_with("}") {
		// FORM A JSON RESPONSE
	}


	// Find user
	// mut user, chk := authorize_user(username, password)

	// mut socket_client := new_client(mut c, 
	// m.clients << socket_client
}

/*
	A sessionID must be generated by authenicating via API Auth Endpoint
*/
pub fn (mut m MessagramServer) client_authenticator(mut c net.TcpConn) 
{
	mut reader := io.new_buffered_reader(reader: c)

	// c.write_string("[ + ] Welcome to Messagram Server v0.0.1\n") or { 0 }
	login := reader.read_line() or { "" }

	println(login)
	if !login.starts_with("{") && !login.ends_with("}") {
		println("[ X ] Error, Invalid login data provided....!\r\n\t=> Disconnecting user " + c.peer_ip() or { "" } + "\r\n\t=>\r\n${login}")
		c.close() or { return }
		return 
	}

	/*
		{
			"cmd_t": ""
			"username": "",
			"sid": "",
			"hwid": "",
			"client_name": "",
			"client_version": ""
		}
	*/
	mut login_data := (jsn.raw_decode("${login}") or { jsn.Any{} }).as_map()

	if "cmd_t" !in login_data || "username" !in login_data || "sid" !in login_data || "hwid" !in login_data {
		println("[ X ] Error, Invalid JSON Response")
		c.close() or { return }
		return
	}

	cmd 		:= (login_data['cmd_t'] 			or { "" }).str()
	username 	:= (login_data['username'] 			or { "" }).str()
	sid 		:= (login_data['sid'] 				or { "" }).str()
	hwid		:= (login_data['hwid'] 				or { "" }).str()
	client_name := (login_data['client_name']		or { "" }).str()
	client_v 	:= (login_data['client_version'] 	or { "" }).str()
	host_addr	:= c.peer_ip() or { "" }

	// Login Authenication
	mut user 		:= m.find_account(username)
	mut client, chk := m.find_client_id(sid, hwid)

	if !chk {
		c.write_string("{\"status\": \"false\", \"resp_t\": \"user_resp\", \"cmd_t\": \"INVALID_LOGIN_INFO\"}") or { 0 }
		c.close() or { return }
		return
	}

	/* Updating the Client's Socket && Client Information */
	m.update_client_info(mut client, mut c, client_name, client_v, mut user)

	mut r := parse_cmd(mut client.info, login)
	mut new_resp := r.parse_cmd_data()

	println("Client Connected ${client}")

	c.write_string("{\"status\": \"true\", \"resp_t\": \"user_resp\", \"cmd_t\": \"SUCCESSFUL_LOGIN\"}") or { 0 }
	m.command_handler(mut c, mut client)
}

/*
	Client Cmd Handler

	Handling account actions such as setting editing, dm actions etc
*/
pub fn (mut m MessagramServer) command_handler(mut socket net.TcpConn, mut client Client)
{
	mut reader := io.new_buffered_reader(reader: socket)
	for
	{
		new_data := reader.read_line() or {
			println("[ X ] Error, Client disconnected from socket\r\n\t=>${client.info.username}.....!")
			m.disconnect_user(mut client.socket)
			return
		}

		println(new_data)
		if !new_data.starts_with("{") || !new_data.ends_with("}")
		{
			println("[ X ] Error, Invalid JSON Data Received!")
			m.disconnect_user(mut client.socket)
			return
		}

		/*
			Default JSON Fields

			There will be additional keys to parse depending on the
			type of commands received
			{
				"cmd": "",
				"username": "",
				"sessionID": "",
				"hwid": "",
				"client_name": "",
				"client_version": ""
			}

			Validate the information below to check the connection
		*/
		json_data 	:= (jsn.raw_decode(new_data) 	or { jsn.Any{} }).as_map()
		cmd 		:= (json_data['cmd_t'] 			or { "" }).str()
		username 	:= (json_data['username'] 		or { "" }).str()
		sid 		:= (json_data['sessionID'] 		or { "" }).str()
		hwid 		:= (json_data['hwid'] 			or { "" }).str() 
		client_name	:= (json_data['client_name']	or { "" }).str()
		client_v	:= (json_data['client_v']		or { "" }).str() 

		// DO ALL CONNECTION VALIDATION CHECKS HERE

		mut r := parse_cmd(mut client.info, new_data)
		mut new_r := r.parse_cmd_data()

		if r.cmd_t == .send_dm_msg { 
			chk := m.send_msg_to_user(mut client, (json_data['to_username'] or { "" }).str(), (json_data['data'] or { "" }).str()) 
			socket.write_string("{\"status\": \"true\", \"resp_t\": \"push_event\", \"cmd_t\": \"send_dm_msg\", \"from_username\": \"Jeff\", \"to_username\": \"vibe\", \"data\": \"gg\"}\n") or { 0 }
			if !chk { 
				println("ERROR: MESSAGE DIDNT SEND")
			}
		}

		println("\x1b[32mOutbound Command: ${m.clients} OUTBOUND END\x1b[39m")

		
		m.clients[0].socket.write_string("gfg\n") or { 0 }

		/* UNCOMMENT THE FUNCTION BELOW ONCE ALL RESPONSES ARE FINISHED */
		
		// handle_command(mut socket, mut new_r)
		// socket.write_string("${new_r.to_str()}") or { 0 }
	}
}

pub fn (mut m MessagramServer) send_msg_to_user(mut from_client Client, to_username string, data string) bool
{
	mut c := 0
	for mut client in m.clients 
	{
		if client.info.username == to_username { 
			println("[ + ] Message Sent to ${to_username} ${client}\nCommand Being Sent: {\"status\": \"true\", \"resp_t\": \"push_event\", \"cmd_t\": \"send_dm_msg\", \"from_username\": \"Jeff\", \"to_username\": \"vibe\", \"data\": \"${data}\"}\n")
			m.clients[c].socket.write_string("{\"status\": \"true\", \"resp_t\": \"push_event\", \"cmd_t\": \"send_dm_msg\", \"from_username\": \"Jeff\", \"to_username\": \"vibe\", \"data\": \"${data}\"}\n")	 or { 0 }
			return true
		}
		c++
	}

	print("failed to send")
	return false
}

pub fn (mut m MessagramServer) disconnect_user(mut socket net.TcpConn) bool
{
	socket.close() or { return false }

	for i, client in m.clients 
	{
		if client.socket == socket { m.clients.delete(i) }
	}

	return true
}

/*
	Find the client id in the (CONNECTED SOCKET CLIENTS) using sid

	Args:
		- sid: sessionID
	
	Returns:
		- Client structure
*/
pub fn (mut m MessagramServer) find_client_id(sid string, h string) (Client, bool)
{
	mut new := Client{socket: &net.TcpConn{}}
	for mut client in m.clients 
	{
		if client.sid == sid && client.hwid == h { return client, true }
	}

	return new, false
}

pub fn (mut m MessagramServer) update_client_info(mut client Client, mut c net.TcpConn, client_name string, client_v string, mut user db.User) 
{
	for mut clnt in m.clients {
		if client.info.username == user.username { 
			clnt.socket 		= c
			clnt.using_app 		= true
			clnt.app_name 		= client_name
			clnt.app_version 	= client_v
			clnt.info 			= user
		}
	}
}

/* 
	Find an account within Messagram's Database (NOT CONNECTED SOCKET CLIENTS)
	
	Args:
		- username: string
	
	Returns:
		- User structure
*/
pub fn (mut m MessagramServer) find_account(username string) db.User
{
	println("Searching... ${username}")
	for mut user in m.users
	{
		if "${user.username}" == "${username}".trim_space() { return user }
	}

	return db.User{}
}