module server

import net

/*
	Handle all commands here. 

	Argument: r has all the JSON data
*/
pub fn handle_command(mut socket net.TcpConn, mut r Response)
{
	// match r.cmd_t
	// {

	// }
}